`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/07/06 15:13:29
// Design Name: 
// Module Name: clz
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module clz(
    input [31:0]a,
    input opt,
    output [31:0] b
    );
  assign b =a[31]==1? 32'h00000000:a[30]==1? 32'h00000001:a[29]==1? 32'h00000002:a[28]==1? 32'h00000003:a[27]==1? 32'h00000004:
            a[26]==1? 32'h00000005:a[25]==1? 32'h00000006:a[24]==1? 32'h00000007:a[23]==1? 32'h00000008:a[22]==1? 32'h00000009:
            a[21]==1? 32'h0000000a:a[20]==1? 32'h0000000b:a[19]==1? 32'h0000000c:a[18]==1? 32'h0000000d:a[17]==1? 32'h0000000e:
            a[16]==1? 32'h0000000f:a[15]==1? 32'h00000010:a[14]==1? 32'h00000011:a[13]==1? 32'h00000012:a[12]==1? 32'h00000013:
            a[11]==1? 32'h00000014:a[10]==1? 32'h00000015:a[9]==1? 32'h00000016:a[8]==1? 32'h00000017:a[7]==1? 32'h00000018:
            a[6]==1? 32'h00000019:a[5]==1? 32'h0000001a:a[4]==1? 32'h0000001b:a[3]==1? 32'h0000001c:a[2]==1? 32'h0000001d:
            a[1]==1? 32'h0000001e:a[0]==1? 32'h0000001f:32'h00000020;
endmodule
